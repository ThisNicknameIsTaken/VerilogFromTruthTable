module DKNF_8_5(i_x0, i_x1, i_x2, i_x3, i_x4, i_x5, i_x6, i_x7, o_y0, o_y1, o_y2, o_y3, o_y4);
	input i_x0, i_x1, i_x2, i_x3, i_x4, i_x5, i_x6, i_x7;
	output o_y0, o_y1, o_y2, o_y3, o_y4;
assign o_y0 = (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7);
assign o_y1 = (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7);
assign o_y2 = (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7);
assign o_y3 = (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7);
assign o_y4 = (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7);
endmodule
