module DDNF_13_8(i_x0, i_x1, i_x2, i_x3, i_x4, i_x5, i_x6, i_x7, i_x8, i_x9, i_x10, i_x11, i_x12, o_y0, o_y1, o_y2, o_y3, o_y4, o_y5, o_y6, o_y7);
	input i_x0, i_x1, i_x2, i_x3, i_x4, i_x5, i_x6, i_x7, i_x8, i_x9, i_x10, i_x11, i_x12;
	output o_y0, o_y1, o_y2, o_y3, o_y4, o_y5, o_y6, o_y7;
assign o_y0 = (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12);
assign o_y1 = (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12);
assign o_y2 = (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12);
assign o_y3 = (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12);
assign o_y4 = (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12);
assign o_y5 = (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12);
assign o_y6 = (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12);
assign o_y7 = (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12) & (~i_x0 | ~i_x1 | ~i_x2 | ~i_x3 | ~i_x4 | ~i_x5 | ~i_x6 | ~i_x7 | ~i_x8 | ~i_x9 | ~i_x10 | ~i_x11 | ~i_x12);
endmodule
